FD-REPOv1	Build time: 1645361143	Applikationer	1
fdimples	0.11.5	FreeDOS installationsprogram - min programvara f�r paketlistredigering	592db6ed
