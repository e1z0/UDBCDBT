Begin3
Language:    SV, 850
Title:       UNFORMAT
Description: Unformat kan �terst�lla en disk som du formaterat av misstag.
Keywords:    format, unformat, h�rddisk,
End
