Begin3
Language:    SV, 850
Title:       more
Description: Visar inneh�llet i en textfil en sida �t g�ngen
Keywords:    freedos, more, sidviare
End
