FD-REPOv1	Build time: 1645361143	Verktyg	5
ambread	20201223	l�sare f�r Ancient Machine Book-formatet	3845698b
callver	2007-08-19a	S�tter DOS-versionen under ett programs k�rning.	b1fd312f
cwsdpmi	7a	32-bitars DPI DOS extender designad f�r DJGPP.	68000114
fdnpkg	0.99.7a	N�tverksbaserad pakethanterare	852ca0c0
v8power	22.02.07	En upps�ttning av f�rb�ttringsverktyg f�r kommandofiler f�r DOS som kan tillhandah�lla textgr�nssnitt och andra behandlingsfunktioner (UPX:at)	50f478fc
