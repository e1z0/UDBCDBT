Begin3
Language:    SV, 850
Title:       DiskCopy
Description: Kopiera en disk eller avbildningsfil till en annan
Keywords:    Freedos, disk, diskcopy, kopiera
End
