Begin3
Language:    SV, 850
Title:       fdxms286
Description: Ers�ttnings-drivrutin f�r XMS f�r '286-system eller b�ttre.
Keywords:    freedos, xms, himem
End
