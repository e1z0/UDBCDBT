FD-REPOv1	Build time: 1645361143	Enhetsdrivrutiner	2
shsufdrv	1.02a	SHSUFDRV �r en drivrutin f�r diskett- och h�rddiskavbildningar. SHSURDRV kopierar avbildningen till RAM och/eller skapar RAM-enheter.	d62292b1
udvd2	2015-03-05d	CD/DVD UltraDMA-enhetsdrivrutin	f17eefb5
