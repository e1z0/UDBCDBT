Begin3
Language:    SV, 850
Title:       devload
Description: Inl�sningprogram f�r drivrutiner p� kommandoraden, har st�d f�r UMB:er
Keywords:    kommandorad, enhet, drivrutin, l�s in, ctload, devload
End
