Begin3
Language:    SV, 850
Title:       Undelete
Description: Undelete l�ter dig �terst�lla borttagna (men �terst�llbara) filer fr�n FAT16/FAT32-filsystem.
Keywords:    undelete, unerase, �terst�ll
End
