Begin3
Language:    SV, 850
Title:       FreeDOS Edit
Description: FreeDOS f�rb�ttrad klon av MS-DOS Edit
Keywords:    redigera, redigerare
End
