Begin3
Language:    SV, 850
Title:       find
Description: Visa alla rader i en eller flera filer som inneh�ller en given str�ng. Omv�nda och skiftl�gesok�nsliga s�kningar ocks� m�jliga.
Keywords:    freedos, hitta, grep
End
