Begin3
Language:    SV, 850
Title:       FreeDOS-k�rnan
Description: FreeDOS-k�rnan
Summary:     FreeDOS-k�rnan (har st�d f�r FAT12/FAT16/FAT32). Inkluderar COUNTRY.SYS, SETVER.SYS och SYS.COM.
Keywords:    k�rna, FreeDOS, DOS, MSDOS
End
