Begin3
Language:    SV, 850
Title:       fc
Description: Filj�mf�relseverktyg
Keywords:    freedos, fil, j�mf�relse, fc
End
