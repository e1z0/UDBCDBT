Begin3
Language:    SV, 850
Title:       attrib
Description: Visa och s�tt filattribut
Keywords:    freedos, attrib
End
