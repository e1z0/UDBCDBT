Begin3
Language:    SV, 850
Title:       swsubst
Description: SUBST och JOIN
Keywords:    freedos, subst, join
End
