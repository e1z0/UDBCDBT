FD-REPOv1	Build time: 1645361143	Arkivprogram	2
unzip	6.00a	Ett fildekomprimeringsverktyg i stil med PKUNZIP.	0a8a4d72
zip	3.0	Ett filarkivprogram i stil med PKZIP.	7efefc96
