Begin3
Language:    SV, 850
Title:       MKEYB
Description: V�ldigt liten tangentbordsdrivrutin, 500-700 byte resident
Keywords:    freedos tangentbord
End
