Begin3
Language:    SV, 850
Title:       Nansi
Description: En ANSI-drivrutin f�r DOS
Keywords:    freedos, nansi, ansi
End
