{

FDIMPLES Language Translation File

Note -- English translations are also built-in to the program. This file is not
required at runtime. However if it is present, settings in here will override
their built-in values.

}

0:SV
1:ogiltig parameter
2:V�nligen v�nta...
3:V�nta
4:Tryck p� en tangent...
5:Grupp
6:Paketmedia hittas ej!
7:Endast installerade paket visas.
8:kan inte hitta pakethanterare FDINST.
9:milj�variabel TEMP �r inte satt.
10:ok�nt
11:installerat
12:Ingen information
13:L�ST
14:Paket
15:inte hittat under
16:V�ntande paketf�r�ndringar:
17:ta bort
18:installera
19:Inga �ndringar.

{ Plural String Values }
20:�ndringar
21:�ndring
22:byte
23:byte
24:Kbyte
25:Kbyte
26:Mbyte
27:Mbyte
28:filer
29:fil
30:k�llkodsfiler
31:k�llkodsfil

{ Basic Load and save stuff }
32:Inkludera paketborttagningar.
33:L�s in anpassningar av paketlista:
34:Spara anpassningar av paketlista:

{ Buttons }
35:OK
36:Avbryt

{ More Status Bar Text }
39:Titel
38:version
39:anv�ndning:
40:[flaggor]

{ Help Messages and such }
50:Publicerat under GNU General Public License, Version 2.0
51:Copyright 2016-2022 Jerome Shidel
52:FDIMPLES tillhandah�ller ett l�ttanv�nt textgr�nssnitt f�r kommandoradspakethanteraren FDINST.

53:Visa denna hj�lpsk�rm.
54:Visa fillista i paketbeskrivning.
55:V�lj att [INTE] automatiskt uppdatera paket.
56:Skapa filer med paketlista f�r anv�ndning med FDI-byggverktyg.
57:Konfigurera FDI installerare BAS och ALLA paketlistor.

58:Tangentbordskommandon f�r anv�ndargr�nssnitt:
59:V�xla markering.
60:�ndra vilket avsnitt eller knapp som har fokus.
61:Flytta fokus ett objekt upp eller ner, �ven Sida upp/ner.
62:Avsluta utan att genomf�r eller spara �ndringar.
63:Visa denna hj�lpsk�rm.
64:V�xla status f�r alla uppdaterbara paket i grupp.
65:V�xla status f�r alla uppdaterbara paket.
66:Visa v�ntade �ndringar.
67:Rensa alla v�ntade �ndringar.
68:Skriv en anpassad paketlistfil som inneh�ller �ndringar.
69:L�s en anpassad paketlistfil och applicera �ndringar.
70:L�t CPU:n sova n�r inget g�rs..
71:Ange enhet eller s�kv�g att anv�nda som arkivk�lla.

{ Package ID's Are all 100 }
100:=Installerat!
100:BASE=FreeDOS Bas
100:ARCHIVER=Arkivprogram
100:BOOT=Uppstartsverktyg
100:DEVEL=Utveckling
100:EDIT=Textredigerare
100:EMULATOR=Emulatorer
100:GAMES=Spel
100:GUI=Grafiska skrivbord
100:NET=N�tverk
100:SOUND=Ljudverktyg
100:UNIXLIKE=Unix-liknande verktyg
100:UTIL=Verktyg
100:UNIX=Unix-liknande verktyg
100:OBSOLETE=F�r�ldrade paket
100:APPS=Applikationer
100:DRIVERS=Enhetsdrivrutiner
