Begin3
Language:    SV, 850
Title:       exe2bin
Description: Konvertera en exe-fil till bin-format
Keywords:    freedos
End
