Begin3
Language:    SV, 850
Title:       GRAPHICS
Description: Till�t Prtscr att skriva ut grafiksk�rmar. (CGA/EGA/VGA/MCGA p� Postskript, ESC/P Epson 8/24-n�lars- och HP PCL-skrivare)
Keywords:    prtscr grafisk skrivardrivrutin dos
End
