Begin3
Language:    SV, 850
Title:       HIMEMX
Description: HimemX �r en XMS-minneshanterar baserade p� FreeDOS Himem.
Keywords:    XMS, himem, minneshanterare
End
